`timescale 1ns/1ps
module uart_tb;

    reg tb_clk_r;
    reg tb_rst_nr;

endmodule /* uart_tb */
