// MIT License
// 
// Copyright (c) 2022 andylithia
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

// Autogenerated MUX tree
module mux7_pyMUX7 (
    input [128-1:0] A,
    input [7-1:0] S,
    output Y
);
wire [64-1:0] mux_level7/* synthesis keep */;
wire [32-1:0] mux_level6/* synthesis keep */;
wire [16-1:0] mux_level5/* synthesis keep */;
wire [8-1:0] mux_level4/* synthesis keep */;
wire [4-1:0] mux_level3/* synthesis keep */;
wire [2-1:0] mux_level2/* synthesis keep */;
wire mux_level1/* synthesis keep */;
genvar gi;
generate
    for(gi=0;gi<64;gi=gi+1) begin : gen_muxl7
        assign mux_level7[gi] = S[0]?mux_level8[2*gi+1]:mux_level8[2*gi];
    end
    for(gi=0;gi<32;gi=gi+1) begin : gen_muxl6
        assign mux_level6[gi] = S[1]?mux_level7[2*gi+1]:mux_level7[2*gi];
    end
    for(gi=0;gi<16;gi=gi+1) begin : gen_muxl5
        assign mux_level5[gi] = S[2]?mux_level6[2*gi+1]:mux_level6[2*gi];
    end
    for(gi=0;gi<8;gi=gi+1) begin : gen_muxl4
        assign mux_level4[gi] = S[3]?mux_level5[2*gi+1]:mux_level5[2*gi];
    end
    for(gi=0;gi<4;gi=gi+1) begin : gen_muxl3
        assign mux_level3[gi] = S[4]?mux_level4[2*gi+1]:mux_level4[2*gi];
    end
    for(gi=0;gi<2;gi=gi+1) begin : gen_muxl2
        assign mux_level2[gi] = S[5]?mux_level3[2*gi+1]:mux_level3[2*gi];
    end
endgenerate
assign mux_level1 = S[6]?mux_level2[1]:mux_level2[0];
assign mux_level7 = A;
assign Y = mux_level1;
endmodule /* mux7_pyMUX7 */